module cpu(
	
);

endmodule