module PraticaV(SW);
	input [17:0] SW;
	
endmodule